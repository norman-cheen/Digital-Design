library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common_pack.all;

ENTITY commandProc IS 
PORT (
    clk:		in std_logic;
    reset:		in std_logic;
    rxNow:		in std_logic;     -- valid (dataReady) signal from Rx
    rxData:			in std_logic_vector (7 downto 0);
    rxDone:		out std_logic;
    numWords_bcd : out BCD_ARRAY_TYPE(2 downto 0); -- bcd output
    aNNN_valid : out std_logic;
    dataReady: in std_logic
    );     
END commandProc;

ARCHITECTURE ANNN of commandProc IS  

  COMPONENT UART_RX_CTRL IS
      PORT(
        RxD: in std_logic;                -- serial data in
        sysclk: in std_logic; 		-- system clock
        reset: in std_logic;		--	synchronous reset
        rxDone: in std_logic;		-- data succesfully read (active high)
        rcvDataReg: out std_logic_vector(7 downto 0); -- received data
        dataReady: out std_logic;	        -- data ready to be read (valid)
        setOE: out std_logic;		-- overrun error (active high)
        setFE: out std_logic		-- frame error (active high)
      );
    END COMPONENT;

    TYPE state_type IS (IDLE, READ_A_a, READ_N1, READ_N2, READ_N3, done1, done2, done3,send_valid);
    SIGNAL curState, nextState: state_type; 
    SIGNAL sig_rxDone, sig_rxNow, sig_ovErr, sig_framErr: std_logic;
    SIGNAL sig_rx: std_logic; 
    SIGNAL sig_rxData: std_logic_vector(7 downto 0);
    SIGNAL bcd_array : BCD_ARRAY_TYPE(2 downto 0);
    
BEGIN
    
  ctrl_nextState: PROCESS(curState, rxData, rxNow)
  BEGIN  
    aNNN_valid <= '0';
    rxDone <= '0';
    
    CASE curState IS 
      
      WHEN IDLE =>
        bcd_array <= ("1111", "1111", "1111");  -- initialise the array
        numWords_bcd <= BCD_array;
        IF rxNow = '1' THEN
          rxDone<= '1';
          IF rxData = X"61" OR rxData = X"41" THEN --in decimal 97(a) and 65(A)
            nextState <= READ_A_a;
          ELSE
            nextState <= IDLE;
          END IF;
        END IF;
        
      WHEN READ_A_a =>
        IF rxNow = '1' THEN
          rxDone<= '1';
          IF ((rxData >= X"30") OR (rxData <= X"39")) THEN
            nextState <= READ_N1;
          ELSIF (rxData = X"61" OR rxData = X"41") THEN
            nextState <= READ_A_a;
          ELSE
            nextState <= IDLE;
          END IF;
        END IF;
      
      WHEN READ_N1 =>
        IF ((rxData = X"30") OR (rxData <= X"39")) THEN
          BCD_array(2) <= rxData(3 downto 0);
          nextState <= done1;
        ELSIF (rxData = X"61" OR rxData = X"41") THEN
          nextState <= READ_A_a;
        ELSE
          nextState <= IDLE;
        END IF;
        
      WHEN done1 => 
        IF rxNow = '1' THEN
          rxDone <= '1';
          nextState <= READ_N2;
        END IF;
      
      WHEN READ_N2 =>
        IF ((rxData = X"30") or (rxData <= X"39")) THEN
          bcd_array(1) <= rxData(3 downto 0);
          nextState <= done2;
        ELSIF rxData = X"61" or rxData = X"41" THEN
          BCD_array(2) <= "1111";
          nextState <= READ_A_a;
        ELSE
          nextState <= IDLE;
        END IF;
        
      WHEN done2 => 
        IF rxNow = '1' THEN
          rxDone <= '1';
          nextState <= READ_N3;
        END IF;
      
      WHEN READ_N3 =>
        IF rxNow = '1' THEN
          IF ((rxData = X"30") or (rxData <= X"39")) THEN
            bcd_array(0) <= rxData(3 downto 0);
            nextState <= done3;
          ELSIF rxData = X"61" or rxData = X"41" THEN
            BCD_array(1) <= "1111";
            BCD_array(2) <= "1111";
            nextState <= READ_A_a;
          ELSE
            nextState <= IDLE;
          END IF;
        END IF;
        
      WHEN done3 => 
        numWords_BCD <= BCD_array;
        rxDone <= '1';
        nextState <= send_valid;
      
      WHEN send_valid =>
        aNNN_valid <= '1';      -- signalling the Nibble Counter to send 'space' after a valid command 
        nextState <= IDLE;

      WHEN OTHERS => 
        nextState <= IDLE;
    END CASE;
  END PROCESS;
  
  stateReg: PROCESS(reset,clk)
  BEGIN
    IF reset = '1'  THEN
      curState <= IDLE;
    ELSIF clk'event AND clk = '1' THEN
      curState <= nextState;
    END IF;
  END PROCESS;

END;   


